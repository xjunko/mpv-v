module main

import gg

const (
	key_toggle_play = [gg.KeyCode.p, gg.KeyCode.space] // not sure, tried to | the enum but v doesnt support it ?
	key_quit        = [gg.KeyCode.q, gg.KeyCode.escape]
)
